library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity divisor_2 is
port(clk:     in     std_logic;
     nRst:    in     std_logic;
     f_out_1: buffer std_logic;
     f_out_2: buffer std_logic);
end entity;

architecture rtl of divisor_2 is
  -- Se�ales
  
begin
  -- Contador modulo 4 con salida de fin de cuenta
  
  
  
  -- Contador m�dulo 3 con entrada de habilitaci�n y salida
  -- de fin de cuenta (independiente de la entrada de habilitaci�n)
   
  
            
end rtl;