-- Autor: TBC
-- Fecha: TBC
-- TBC
-- TBC

library ieee;
use ieee.std_logic_1164.all;

entity reg16b_ena_rst is
port(
  clk : TBC;
  nRST: TBC;
  sRST: TBC;
  ena : TBC;
  Din : TBC;
  Dout: TBC
);
end entity;

architecture TBC of TBC is
begin

   process(TBC)
   begin
      if TBC
	     TBC
      elsif TBC then
         if TBC then
           Dout <=(others => '0');
         elsif TBC then
           Dout <= Din;
         end if;
      end if;
   end process;
end rtl;